��/ *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ i n _ r o u t e r _ 0 _ o u t 0 ;  
 w i r e   c b _ i n _ r o u t e r _ 0 _ o u t 1 ;  
 w i r e   c b _ i n _ r o u t e r _ 0 _ o u t 2 ;  
 w i r e   c b _ i n _ r o u t e r _ 0 _ o u t 3 ;  
 w i r e   [ 0 : 5 ]   c b _ i n _ r o u t e r _ 0 _ s e l ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ o u t _ r o u t e r _ 0 _ i n 0 ;  
 w i r e   c b _ o u t _ r o u t e r _ 0 _ i n 1 ;  
 w i r e   c b _ o u t _ r o u t e r _ 0 _ i n 2 ;  
 w i r e   c b _ o u t _ r o u t e r _ 0 _ i n 3 ;  
 w i r e   [ 0 : 5 ]   c b _ o u t _ r o u t e r _ 0 _ s e l ;  
  
  
 D e m o 1 _ a l t e r a _ m e r l i n _ r o u t e r _ 1 9 2 0 _ e n 6 j v e a   r o u t e r _ 0 0 1   (  
 	   . s i n k _ v a l i d ( c b _ i n _ r o u t e r _ 0 _ o u t 0 ) ,  
 	   . s i n k _ s t a r t o f p a c k e t ( c b _ i n _ r o u t e r _ 0 _ o u t 1 ) ,  
 	   . s i n k _ e n d o f p a c k e t ( c b _ i n _ r o u t e r _ 0 _ o u t 2 ) ,  
 	   . s r c _ r e a d y ( c b _ i n _ r o u t e r _ 0 _ o u t 3 ) ,  
 	   . s i n k _ r e a d y ( c b _ o u t _ r o u t e r _ 0 _ i n 0 ) ,  
 	   . s r c _ v a l i d ( c b _ o u t _ r o u t e r _ 0 _ i n 1 ) ,  
 	   . s r c _ s t a r t o f p a c k e t ( c b _ o u t _ r o u t e r _ 0 _ i n 2 ) ,  
 	   . s r c _ e n d o f p a c k e t ( c b _ o u t _ r o u t e r _ 0 _ i n 3 ) ,  
 	   . s i n k _ d a t a ( i n t e l _ n i o s v _ m _ 0 _ d a t a _ m a n a g e r _ a g e n t _ r e a d _ c p _ d a t a ) ,  
 	   . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	   . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	   . s r c _ d a t a ( r o u t e r _ 0 0 1 _ s r c _ d a t a ) ,  
 	   . s r c _ c h a n n e l ( r o u t e r _ 0 0 1 _ s r c _ c h a n n e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ i n _ r o u t e r _ 0   (  
 	   . i n 0 ( i n t e l _ n i o s v _ m _ 0 _ d a t a _ m a n a g e r _ a g e n t _ r e a d _ c p _ s t a r t o f p a c k e t ) ,  
 	   . i n 1 ( i n t e l _ n i o s v _ m _ 0 _ d a t a _ m a n a g e r _ a g e n t _ r e a d _ c p _ e n d o f p a c k e t ) ,  
 	   . i n 2 ( r o u t e r _ 0 0 1 _ s r c _ r e a d y ) ,  
 	   . i n 3 ( i n t e l _ n i o s v _ m _ 0 _ d a t a _ m a n a g e r _ a g e n t _ r e a d _ c p _ v a l i d ) ,  
 	   . o u t 0 ( c b _ i n _ r o u t e r _ 0 _ o u t 0 ) ,  
 	   . o u t 1 ( c b _ i n _ r o u t e r _ 0 _ o u t 1 ) ,  
 	   . o u t 2 ( c b _ i n _ r o u t e r _ 0 _ o u t 2 ) ,  
 	   . o u t 3 ( c b _ i n _ r o u t e r _ 0 _ o u t 3 ) ,  
 	   . s e l 0 ( c b _ i n _ r o u t e r _ 0 _ s e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ o u t _ r o u t e r _ 0   (  
 	   . i n 0 ( c b _ o u t _ r o u t e r _ 0 _ i n 0 ) ,  
 	   . i n 1 ( c b _ o u t _ r o u t e r _ 0 _ i n 1 ) ,  
 	   . i n 2 ( c b _ o u t _ r o u t e r _ 0 _ i n 2 ) ,  
 	   . i n 3 ( c b _ o u t _ r o u t e r _ 0 _ i n 3 ) ,  
 	   . o u t 0 ( s i n k _ r e a d y ) ,  
 	   . o u t 1 ( s r c _ v a l i d ) ,  
 	   . o u t 2 ( s r c _ s t a r t o f p a c k e t ) ,  
 	   . o u t 3 ( s r c _ e n d o f p a c k e t ) ,  
 	   . s e l 0 ( c b _ o u t _ r o u t e r _ 0 _ s e l )  
 ) ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ i n _ r o u t e r _ 1 _ o u t 0 ;  
 w i r e   c b _ i n _ r o u t e r _ 1 _ o u t 1 ;  
 w i r e   c b _ i n _ r o u t e r _ 1 _ o u t 2 ;  
 w i r e   c b _ i n _ r o u t e r _ 1 _ o u t 3 ;  
 w i r e   [ 0 : 5 ]   c b _ i n _ r o u t e r _ 1 _ s e l ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ o u t _ r o u t e r _ 1 _ i n 0 ;  
 w i r e   c b _ o u t _ r o u t e r _ 1 _ i n 1 ;  
 w i r e   c b _ o u t _ r o u t e r _ 1 _ i n 2 ;  
 w i r e   c b _ o u t _ r o u t e r _ 1 _ i n 3 ;  
 w i r e   [ 0 : 5 ]   c b _ o u t _ r o u t e r _ 1 _ s e l ;  
  
  
 D e m o 1 _ a l t e r a _ m e r l i n _ r o u t e r _ 1 9 2 0 _ k x o v a a y   r o u t e r _ 0 0 2   (  
 	   . s i n k _ v a l i d ( c b _ i n _ r o u t e r _ 1 _ o u t 0 ) ,  
 	   . s i n k _ s t a r t o f p a c k e t ( c b _ i n _ r o u t e r _ 1 _ o u t 1 ) ,  
 	   . s i n k _ e n d o f p a c k e t ( c b _ i n _ r o u t e r _ 1 _ o u t 2 ) ,  
 	   . s r c _ r e a d y ( c b _ i n _ r o u t e r _ 1 _ o u t 3 ) ,  
 	   . s i n k _ r e a d y ( c b _ o u t _ r o u t e r _ 1 _ i n 0 ) ,  
 	   . s r c _ v a l i d ( c b _ o u t _ r o u t e r _ 1 _ i n 1 ) ,  
 	   . s r c _ s t a r t o f p a c k e t ( c b _ o u t _ r o u t e r _ 1 _ i n 2 ) ,  
 	   . s r c _ e n d o f p a c k e t ( c b _ o u t _ r o u t e r _ 1 _ i n 3 ) ,  
 	   . s i n k _ d a t a ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ w r i t e _ c p _ d a t a ) ,  
 	   . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	   . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	   . s r c _ d a t a ( r o u t e r _ 0 0 2 _ s r c _ d a t a ) ,  
 	   . s r c _ c h a n n e l ( r o u t e r _ 0 0 2 _ s r c _ c h a n n e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ i n _ r o u t e r _ 1   (  
 	   . i n 0 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ w r i t e _ c p _ s t a r t o f p a c k e t ) ,  
 	   . i n 1 ( r o u t e r _ 0 0 2 _ s r c _ r e a d y ) ,  
 	   . i n 2 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ w r i t e _ c p _ e n d o f p a c k e t ) ,  
 	   . i n 3 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ w r i t e _ c p _ v a l i d ) ,  
 	   . o u t 0 ( c b _ i n _ r o u t e r _ 1 _ o u t 0 ) ,  
 	   . o u t 1 ( c b _ i n _ r o u t e r _ 1 _ o u t 1 ) ,  
 	   . o u t 2 ( c b _ i n _ r o u t e r _ 1 _ o u t 2 ) ,  
 	   . o u t 3 ( c b _ i n _ r o u t e r _ 1 _ o u t 3 ) ,  
 	   . s e l 0 ( c b _ i n _ r o u t e r _ 1 _ s e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ o u t _ r o u t e r _ 1   (  
 	   . i n 0 ( c b _ o u t _ r o u t e r _ 1 _ i n 0 ) ,  
 	   . i n 1 ( c b _ o u t _ r o u t e r _ 1 _ i n 1 ) ,  
 	   . i n 2 ( c b _ o u t _ r o u t e r _ 1 _ i n 2 ) ,  
 	   . i n 3 ( c b _ o u t _ r o u t e r _ 1 _ i n 3 ) ,  
 	   . o u t 0 ( s i n k _ r e a d y ) ,  
 	   . o u t 1 ( s r c _ v a l i d ) ,  
 	   . o u t 2 ( s r c _ s t a r t o f p a c k e t ) ,  
 	   . o u t 3 ( s r c _ e n d o f p a c k e t ) ,  
 	   . s e l 0 ( c b _ o u t _ r o u t e r _ 1 _ s e l )  
 ) ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ i n _ r o u t e r _ 2 _ o u t 0 ;  
 w i r e   c b _ i n _ r o u t e r _ 2 _ o u t 1 ;  
 w i r e   c b _ i n _ r o u t e r _ 2 _ o u t 2 ;  
 w i r e   c b _ i n _ r o u t e r _ 2 _ o u t 3 ;  
 w i r e   [ 0 : 5 ]   c b _ i n _ r o u t e r _ 2 _ s e l ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ o u t _ r o u t e r _ 2 _ i n 0 ;  
 w i r e   c b _ o u t _ r o u t e r _ 2 _ i n 1 ;  
 w i r e   c b _ o u t _ r o u t e r _ 2 _ i n 2 ;  
 w i r e   c b _ o u t _ r o u t e r _ 2 _ i n 3 ;  
 w i r e   [ 0 : 5 ]   c b _ o u t _ r o u t e r _ 2 _ s e l ;  
  
  
 D e m o 1 _ a l t e r a _ m e r l i n _ r o u t e r _ 1 9 2 0 _ k x o v a a y   r o u t e r _ 0 0 3   (  
 	   . s i n k _ v a l i d ( c b _ i n _ r o u t e r _ 2 _ o u t 0 ) ,  
 	   . s i n k _ s t a r t o f p a c k e t ( c b _ i n _ r o u t e r _ 2 _ o u t 1 ) ,  
 	   . s i n k _ e n d o f p a c k e t ( c b _ i n _ r o u t e r _ 2 _ o u t 2 ) ,  
 	   . s r c _ r e a d y ( c b _ i n _ r o u t e r _ 2 _ o u t 3 ) ,  
 	   . s i n k _ r e a d y ( c b _ o u t _ r o u t e r _ 2 _ i n 0 ) ,  
 	   . s r c _ v a l i d ( c b _ o u t _ r o u t e r _ 2 _ i n 1 ) ,  
 	   . s r c _ s t a r t o f p a c k e t ( c b _ o u t _ r o u t e r _ 2 _ i n 2 ) ,  
 	   . s r c _ e n d o f p a c k e t ( c b _ o u t _ r o u t e r _ 2 _ i n 3 ) ,  
 	   . s i n k _ d a t a ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ r e a d _ c p _ d a t a ) ,  
 	   . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	   . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	   . s r c _ d a t a ( r o u t e r _ 0 0 3 _ s r c _ d a t a ) ,  
 	   . s r c _ c h a n n e l ( r o u t e r _ 0 0 3 _ s r c _ c h a n n e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ i n _ r o u t e r _ 2   (  
 	   . i n 0 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ r e a d _ c p _ s t a r t o f p a c k e t ) ,  
 	   . i n 1 ( r o u t e r _ 0 0 3 _ s r c _ r e a d y ) ,  
 	   . i n 2 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ r e a d _ c p _ v a l i d ) ,  
 	   . i n 3 ( i n t e l _ n i o s v _ m _ 0 _ i n s t r u c t i o n _ m a n a g e r _ a g e n t _ r e a d _ c p _ e n d o f p a c k e t ) ,  
 	   . o u t 0 ( c b _ i n _ r o u t e r _ 2 _ o u t 0 ) ,  
 	   . o u t 1 ( c b _ i n _ r o u t e r _ 2 _ o u t 1 ) ,  
 	   . o u t 2 ( c b _ i n _ r o u t e r _ 2 _ o u t 2 ) ,  
 	   . o u t 3 ( c b _ i n _ r o u t e r _ 2 _ o u t 3 ) ,  
 	   . s e l 0 ( c b _ i n _ r o u t e r _ 2 _ s e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ o u t _ r o u t e r _ 2   (  
 	   . i n 0 ( c b _ o u t _ r o u t e r _ 2 _ i n 0 ) ,  
 	   . i n 1 ( c b _ o u t _ r o u t e r _ 2 _ i n 1 ) ,  
 	   . i n 2 ( c b _ o u t _ r o u t e r _ 2 _ i n 2 ) ,  
 	   . i n 3 ( c b _ o u t _ r o u t e r _ 2 _ i n 3 ) ,  
 	   . o u t 0 ( s i n k _ r e a d y ) ,  
 	   . o u t 1 ( s r c _ v a l i d ) ,  
 	   . o u t 2 ( s r c _ s t a r t o f p a c k e t ) ,  
 	   . o u t 3 ( s r c _ e n d o f p a c k e t ) ,  
 	   . s e l 0 ( c b _ o u t _ r o u t e r _ 2 _ s e l )  
 ) ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ i n _ r o u t e r _ 3 _ o u t 0 ;  
 w i r e   c b _ i n _ r o u t e r _ 3 _ o u t 1 ;  
 w i r e   c b _ i n _ r o u t e r _ 3 _ o u t 2 ;  
 w i r e   c b _ i n _ r o u t e r _ 3 _ o u t 3 ;  
 w i r e   [ 0 : 5 ]   c b _ i n _ r o u t e r _ 3 _ s e l ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ o u t _ r o u t e r _ 3 _ i n 0 ;  
 w i r e   c b _ o u t _ r o u t e r _ 3 _ i n 1 ;  
 w i r e   c b _ o u t _ r o u t e r _ 3 _ i n 2 ;  
 w i r e   c b _ o u t _ r o u t e r _ 3 _ i n 3 ;  
 w i r e   [ 0 : 5 ]   c b _ o u t _ r o u t e r _ 3 _ s e l ;  
  
  
 D e m o 1 _ a l t e r a _ m e r l i n _ r o u t e r _ 1 9 2 0 _ 7 i o 6 p 2 i   r o u t e r _ 0 0 7   (  
 	   . s i n k _ v a l i d ( c b _ i n _ r o u t e r _ 3 _ o u t 0 ) ,  
 	   . s i n k _ s t a r t o f p a c k e t ( c b _ i n _ r o u t e r _ 3 _ o u t 1 ) ,  
 	   . s i n k _ e n d o f p a c k e t ( c b _ i n _ r o u t e r _ 3 _ o u t 2 ) ,  
 	   . s r c _ r e a d y ( c b _ i n _ r o u t e r _ 3 _ o u t 3 ) ,  
 	   . s i n k _ r e a d y ( c b _ o u t _ r o u t e r _ 3 _ i n 0 ) ,  
 	   . s r c _ v a l i d ( c b _ o u t _ r o u t e r _ 3 _ i n 1 ) ,  
 	   . s r c _ s t a r t o f p a c k e t ( c b _ o u t _ r o u t e r _ 3 _ i n 2 ) ,  
 	   . s r c _ e n d o f p a c k e t ( c b _ o u t _ r o u t e r _ 3 _ i n 3 ) ,  
 	   . s i n k _ d a t a ( i n t e l _ n i o s v _ m _ 0 _ t i m e r _ s w _ a g e n t _ a g e n t _ r p _ d a t a ) ,  
 	   . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	   . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	   . s r c _ d a t a ( r o u t e r _ 0 0 7 _ s r c _ d a t a ) ,  
 	   . s r c _ c h a n n e l ( r o u t e r _ 0 0 7 _ s r c _ c h a n n e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ i n _ r o u t e r _ 3   (  
 	   . i n 0 ( i n t e l _ n i o s v _ m _ 0 _ t i m e r _ s w _ a g e n t _ a g e n t _ r p _ s t a r t o f p a c k e t ) ,  
 	   . i n 1 ( i n t e l _ n i o s v _ m _ 0 _ t i m e r _ s w _ a g e n t _ a g e n t _ r p _ v a l i d ) ,  
 	   . i n 2 ( i n t e l _ n i o s v _ m _ 0 _ t i m e r _ s w _ a g e n t _ a g e n t _ r p _ e n d o f p a c k e t ) ,  
 	   . i n 3 ( r o u t e r _ 0 0 7 _ s r c _ r e a d y ) ,  
 	   . o u t 0 ( c b _ i n _ r o u t e r _ 3 _ o u t 0 ) ,  
 	   . o u t 1 ( c b _ i n _ r o u t e r _ 3 _ o u t 1 ) ,  
 	   . o u t 2 ( c b _ i n _ r o u t e r _ 3 _ o u t 2 ) ,  
 	   . o u t 3 ( c b _ i n _ r o u t e r _ 3 _ o u t 3 ) ,  
 	   . s e l 0 ( c b _ i n _ r o u t e r _ 3 _ s e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ o u t _ r o u t e r _ 3   (  
 	   . i n 0 ( c b _ o u t _ r o u t e r _ 3 _ i n 0 ) ,  
 	   . i n 1 ( c b _ o u t _ r o u t e r _ 3 _ i n 1 ) ,  
 	   . i n 2 ( c b _ o u t _ r o u t e r _ 3 _ i n 2 ) ,  
 	   . i n 3 ( c b _ o u t _ r o u t e r _ 3 _ i n 3 ) ,  
 	   . o u t 0 ( s i n k _ r e a d y ) ,  
 	   . o u t 1 ( s r c _ v a l i d ) ,  
 	   . o u t 2 ( s r c _ s t a r t o f p a c k e t ) ,  
 	   . o u t 3 ( s r c _ e n d o f p a c k e t ) ,  
 	   . s e l 0 ( c b _ o u t _ r o u t e r _ 3 _ s e l )  
 ) ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ i n _ r o u t e r _ 4 _ o u t 0 ;  
 w i r e   c b _ i n _ r o u t e r _ 4 _ o u t 1 ;  
 w i r e   c b _ i n _ r o u t e r _ 4 _ o u t 2 ;  
 w i r e   c b _ i n _ r o u t e r _ 4 _ o u t 3 ;  
 w i r e   [ 0 : 5 ]   c b _ i n _ r o u t e r _ 4 _ s e l ;  
  
  
 / *   P r i n t i n g   w i r e s           * /  
 w i r e   c b _ o u t _ r o u t e r _ 4 _ i n 0 ;  
 w i r e   c b _ o u t _ r o u t e r _ 4 _ i n 1 ;  
 w i r e   c b _ o u t _ r o u t e r _ 4 _ i n 2 ;  
 w i r e   c b _ o u t _ r o u t e r _ 4 _ i n 3 ;  
 w i r e   [ 0 : 5 ]   c b _ o u t _ r o u t e r _ 4 _ s e l ;  
  
  
 D e m o 1 _ a l t e r a _ m e r l i n _ r o u t e r _ 1 9 2 0 _ 7 i o 6 p 2 i   r o u t e r _ 0 0 4   (  
 	   . s i n k _ v a l i d ( c b _ i n _ r o u t e r _ 4 _ o u t 0 ) ,  
 	   . s i n k _ s t a r t o f p a c k e t ( c b _ i n _ r o u t e r _ 4 _ o u t 1 ) ,  
 	   . s i n k _ e n d o f p a c k e t ( c b _ i n _ r o u t e r _ 4 _ o u t 2 ) ,  
 	   . s r c _ r e a d y ( c b _ i n _ r o u t e r _ 4 _ o u t 3 ) ,  
 	   . s i n k _ r e a d y ( c b _ o u t _ r o u t e r _ 4 _ i n 0 ) ,  
 	   . s r c _ v a l i d ( c b _ o u t _ r o u t e r _ 4 _ i n 1 ) ,  
 	   . s r c _ s t a r t o f p a c k e t ( c b _ o u t _ r o u t e r _ 4 _ i n 2 ) ,  
 	   . s r c _ e n d o f p a c k e t ( c b _ o u t _ r o u t e r _ 4 _ i n 3 ) ,  
 	   . s i n k _ d a t a ( j t a g _ u a r t _ 0 _ a v a l o n _ j t a g _ s l a v e _ a g e n t _ r p _ d a t a ) ,  
 	   . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	   . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	   . s r c _ d a t a ( r o u t e r _ 0 0 4 _ s r c _ d a t a ) ,  
 	   . s r c _ c h a n n e l ( r o u t e r _ 0 0 4 _ s r c _ c h a n n e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ i n _ r o u t e r _ 4   (  
 	   . i n 0 ( j t a g _ u a r t _ 0 _ a v a l o n _ j t a g _ s l a v e _ a g e n t _ r p _ v a l i d ) ,  
 	   . i n 1 ( j t a g _ u a r t _ 0 _ a v a l o n _ j t a g _ s l a v e _ a g e n t _ r p _ e n d o f p a c k e t ) ,  
 	   . i n 2 ( j t a g _ u a r t _ 0 _ a v a l o n _ j t a g _ s l a v e _ a g e n t _ r p _ s t a r t o f p a c k e t ) ,  
 	   . i n 3 ( r o u t e r _ 0 0 4 _ s r c _ r e a d y ) ,  
 	   . o u t 0 ( c b _ i n _ r o u t e r _ 4 _ o u t 0 ) ,  
 	   . o u t 1 ( c b _ i n _ r o u t e r _ 4 _ o u t 1 ) ,  
 	   . o u t 2 ( c b _ i n _ r o u t e r _ 4 _ o u t 2 ) ,  
 	   . o u t 3 ( c b _ i n _ r o u t e r _ 4 _ o u t 3 ) ,  
 	   . s e l 0 ( c b _ i n _ r o u t e r _ 4 _ s e l )  
 ) ;  
  
  
 c r b a r 4 x 4   c b _ o u t _ r o u t e r _ 4   (  
 	   . i n 0 ( c b _ o u t _ r o u t e r _ 4 _ i n 0 ) ,  
 	   . i n 1 ( c b _ o u t _ r o u t e r _ 4 _ i n 1 ) ,  
 	   . i n 2 ( c b _ o u t _ r o u t e r _ 4 _ i n 2 ) ,  
 	   . i n 3 ( c b _ o u t _ r o u t e r _ 4 _ i n 3 ) ,  
 	   . o u t 0 ( s i n k _ r e a d y ) ,  
 	   . o u t 1 ( s r c _ v a l i d ) ,  
 	   . o u t 2 ( s r c _ s t a r t o f p a c k e t ) ,  
 	   . o u t 3 ( s r c _ e n d o f p a c k e t ) ,  
 	   . s e l 0 ( c b _ o u t _ r o u t e r _ 4 _ s e l )  
 ) ;  
  
  
 w i r e   [ 5 9 : 0 ]   s e l e c t _ l i n e s ;  
  
 a s s i g n   c b _ i n _ r o u t e r _ 0 _ s e l   =   s e l e c t _ l i n e s [ 5 : 0 ] ;  
 a s s i g n   c b _ o u t _ r o u t e r _ 0 _ s e l   =   s e l e c t _ l i n e s [ 1 1 : 6 ] ;  
 a s s i g n   c b _ i n _ r o u t e r _ 1 _ s e l   =   s e l e c t _ l i n e s [ 1 7 : 1 2 ] ;  
 a s s i g n   c b _ o u t _ r o u t e r _ 1 _ s e l   =   s e l e c t _ l i n e s [ 2 3 : 1 8 ] ;  
 a s s i g n   c b _ i n _ r o u t e r _ 2 _ s e l   =   s e l e c t _ l i n e s [ 2 9 : 2 4 ] ;  
 a s s i g n   c b _ o u t _ r o u t e r _ 2 _ s e l   =   s e l e c t _ l i n e s [ 3 5 : 3 0 ] ;  
 a s s i g n   c b _ i n _ r o u t e r _ 3 _ s e l   =   s e l e c t _ l i n e s [ 4 1 : 3 6 ] ;  
 a s s i g n   c b _ o u t _ r o u t e r _ 3 _ s e l   =   s e l e c t _ l i n e s [ 4 7 : 4 2 ] ;  
 a s s i g n   c b _ i n _ r o u t e r _ 4 _ s e l   =   s e l e c t _ l i n e s [ 5 3 : 4 8 ] ;  
 a s s i g n   c b _ o u t _ r o u t e r _ 4 _ s e l   =   s e l e c t _ l i n e s [ 5 9 : 5 4 ] ;  
  
 a c t i v a t i o n _ p a c k a g e _ n _ b i t   a c t 1   (  
 	 . c l k ( c l o c k _ i n _ o u t _ c l k _ c l k ) ,  
 	 . r e s e t ( i n t e l _ n i o s v _ m _ 0 _ r e s e t _ r e s e t _ b r i d g e _ i n _ r e s e t _ r e s e t ) ,  
 	 . s e r i a l _ i n ( s e r i a l _ i n ) ,  
 	 . p a r a l l e l _ o u t ( s e l e c t _ l i n e s )  
 ) ;  
 